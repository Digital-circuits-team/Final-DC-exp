module(clk,newCh);
    input clk;
    output [23:0] randomNum;

    


endmodule